// Verilog test fixture created from schematic E:\Adam\GitHubLocallReopsitory\EngineerSoftCPU\APCPU\MainCPU.sch - Sat Jan 16 13:22:42 2021

`timescale 1ns / 1ps

module MainCPU_MainCPU_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   MainCPU UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
